dimensions:
	time = UNLIMITED ; // (10 currently)
	time_0 = 20 ;
variables:
	double temp(time) ;
		temp:standard_name = "air_temperature" ;
		temp:units = "K" ;
	int64 time(time) ;
		time:units = "1" ;
		time:standard_name = "time" ;
	double temp2(time_0) ;
		temp2:long_name = "air_temperature" ;
		temp2:units = "K" ;
	int64 time_0(time_0) ;
		time_0:units = "1" ;
		time_0:standard_name = "time" ;
	double temp3(time) ;
		temp3:long_name = "air_temperature" ;
		temp3:units = "K" ;

// global attributes:
		:Conventions = "CF-1.5" ;
}
